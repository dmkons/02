library ieee;
use ieee.stdd_logic_1164.all;


entity processor is
end processor;

architecture Behavioral of processor is
begin
end Behavioral;

